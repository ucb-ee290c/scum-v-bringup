module SCUMVTuning(
  output        auto_mmio_in_a_ready,
  input         auto_mmio_in_a_valid,
  input  [2:0]  auto_mmio_in_a_bits_opcode,
                auto_mmio_in_a_bits_param,
  input  [1:0]  auto_mmio_in_a_bits_size,
  input  [15:0] auto_mmio_in_a_bits_source,
                auto_mmio_in_a_bits_address,
  input  [3:0]  auto_mmio_in_a_bits_mask,
  input  [31:0] auto_mmio_in_a_bits_data,
  input         auto_mmio_in_a_bits_corrupt,
                auto_mmio_in_d_ready,
  output        auto_mmio_in_d_valid,
  output [2:0]  auto_mmio_in_d_bits_opcode,
  output [1:0]  auto_mmio_in_d_bits_size,
  output [15:0] auto_mmio_in_d_bits_source,
  output [31:0] auto_mmio_in_d_bits_data,
  input         auto_clock_in_clock,
                auto_clock_in_reset,
  output [8:0]  io_oscillator_tuneOut_adc_coarse,	
  output [5:0]  io_oscillator_tuneOut_dig,	
  output [1:0]  io_oscillator_tuneOut_cpuSel,	
  output        io_oscillator_reset_adc,	
                io_oscillator_reset_dig,	
  output [4:0]  io_supply_bgr_tempCtrl,	
                io_supply_bgr_vrefCtrl,	
                io_supply_currentSrc_leftCtrl,	
                io_supply_currentSrc_rightCtrl,	
  output        io_supply_clkOvrd,	
                io_radar_rampGenerator_clkMuxSel,	
                io_radar_rampGenerator_enable,	
  output [7:0]  io_radar_rampGenerator_frequencyStepStart,	
                io_radar_rampGenerator_numFrequencySteps,	
  output [23:0] io_radar_rampGenerator_numCyclesPerFrequency,	
  output [31:0] io_radar_rampGenerator_numIdleCycles,	
  output        io_radar_rampGenerator_rst,	
  output [5:0]  io_radar_rampGenerator_idac_control,	
  output [1:0]  io_radar_rampGenerator_rx_out_sel,	
  output [4:0]  io_radar_vco_capTuning,	
  output        io_radar_vco_enable,	
                io_radar_vco_divEnable,	
                io_radar_pa_enable,	
                io_radar_pa_bypass,	
                io_radar_pa_inputMuxSel,	
                io_radar_clkOvrd	
);

  SCUMVTuningFrontend scumvtuningFrontend (	// @[generators/scumvtuning/src/main/scala/SCUMVTuning.scala:312:39]
    .clock                                        (auto_clock_in_clock),
    .reset                                        (auto_clock_in_reset),
    .auto_control_xing_in_a_ready                 (auto_mmio_in_a_ready),
    .auto_control_xing_in_a_valid                 (auto_mmio_in_a_valid),
    .auto_control_xing_in_a_bits_opcode           (auto_mmio_in_a_bits_opcode),
    .auto_control_xing_in_a_bits_param            (auto_mmio_in_a_bits_param),
    .auto_control_xing_in_a_bits_size             (auto_mmio_in_a_bits_size),
    .auto_control_xing_in_a_bits_source           (auto_mmio_in_a_bits_source),
    .auto_control_xing_in_a_bits_address          (auto_mmio_in_a_bits_address),
    .auto_control_xing_in_a_bits_mask             (auto_mmio_in_a_bits_mask),
    .auto_control_xing_in_a_bits_data             (auto_mmio_in_a_bits_data),
    .auto_control_xing_in_a_bits_corrupt          (auto_mmio_in_a_bits_corrupt),
    .auto_control_xing_in_d_ready                 (auto_mmio_in_d_ready),
    .auto_control_xing_in_d_valid                 (auto_mmio_in_d_valid),
    .auto_control_xing_in_d_bits_opcode           (auto_mmio_in_d_bits_opcode),
    .auto_control_xing_in_d_bits_size             (auto_mmio_in_d_bits_size),
    .auto_control_xing_in_d_bits_source           (auto_mmio_in_d_bits_source),
    .auto_control_xing_in_d_bits_data             (auto_mmio_in_d_bits_data),
    .io_oscillator_tuneOut_adc_coarse             (io_oscillator_tuneOut_adc_coarse),
    .io_oscillator_tuneOut_dig                    (io_oscillator_tuneOut_dig),
    .io_oscillator_tuneOut_cpuSel                 (io_oscillator_tuneOut_cpuSel),
    .io_oscillator_reset_adc                      (io_oscillator_reset_adc),
    .io_oscillator_reset_dig                      (io_oscillator_reset_dig),
    .io_supply_bgr_tempCtrl                       (io_supply_bgr_tempCtrl),
    .io_supply_bgr_vrefCtrl                       (io_supply_bgr_vrefCtrl),
    .io_supply_currentSrc_leftCtrl                (io_supply_currentSrc_leftCtrl),
    .io_supply_currentSrc_rightCtrl               (io_supply_currentSrc_rightCtrl),
    .io_supply_clkOvrd                            (io_supply_clkOvrd),
    .io_radar_rampGenerator_clkMuxSel             (io_radar_rampGenerator_clkMuxSel),
    .io_radar_rampGenerator_enable                (io_radar_rampGenerator_enable),
    .io_radar_rampGenerator_frequencyStepStart    (io_radar_rampGenerator_frequencyStepStart),
    .io_radar_rampGenerator_numFrequencySteps     (io_radar_rampGenerator_numFrequencySteps),
    .io_radar_rampGenerator_numCyclesPerFrequency (io_radar_rampGenerator_numCyclesPerFrequency),
    .io_radar_rampGenerator_numIdleCycles         (io_radar_rampGenerator_numIdleCycles),
    .io_radar_rampGenerator_rst                   (io_radar_rampGenerator_rst),
    .io_radar_rampGenerator_idac_control          (io_radar_rampGenerator_idac_control),
    .io_radar_rampGenerator_rx_out_sel            (io_radar_rampGenerator_rx_out_sel),
    .io_radar_vco_capTuning                       (io_radar_vco_capTuning),
    .io_radar_vco_enable                          (io_radar_vco_enable),
    .io_radar_vco_divEnable                       (io_radar_vco_divEnable),
    .io_radar_pa_enable                           (io_radar_pa_enable),
    .io_radar_pa_bypass                           (io_radar_pa_bypass),
    .io_radar_pa_inputMuxSel                      (io_radar_pa_inputMuxSel),
    .io_radar_clkOvrd                             (io_radar_clkOvrd)
  );
endmodule

