`timescale 1ns / 1ps

// Helper module: Ready/Valid backpressure ready gater with pattern
module rv_ready_gate #(parameter integer PATTERN_LEN = 9) (
    input  wire        clock,
    input  wire        reset,
    input  wire        enable,
    input  wire [8:0]  pattern,
    input  wire        valid_in,
    input  wire        raw_ready_in,
    output reg  [3:0]  index,
    output wire        ready_gated_out
);
    always @(posedge clock) begin
        if (reset) begin
            index <= 4'd0;
        end else if (enable) begin
            // Advance index only when there is an actual transaction attempt (valid & raw ready)
            if (valid_in && raw_ready_in) begin
                if (index >= PATTERN_LEN - 1)
                    index <= 4'd0;
                else
                    index <= index + 1'b1;
            end
        end
    end

    assign ready_gated_out = enable ? (raw_ready_in & pattern[index]) : raw_ready_in;
endmodule

// Helper module: Backpressure counters and event logging
module rv_bp_counters (
    input  wire        clock,
    input  wire        reset,
    input  wire        enable,
    input  wire        valid_in,
    input  wire        raw_ready_in,
    input  wire        ready_gated_in,
    input  integer     tb_log_fd,
    output reg  [31:0] backpressure_events,
    output reg  [31:0] transactions_accepted,
    output reg  [31:0] transactions_stalled
);
    always @(posedge clock) begin
        if (reset) begin
            backpressure_events   <= 32'd0;
            transactions_accepted <= 32'd0;
            transactions_stalled  <= 32'd0;
        end else if (enable) begin
            // Backpressure event when raw ready is high, but gated ready is low while valid is asserted
            if (valid_in && raw_ready_in && !ready_gated_in) begin
                backpressure_events <= backpressure_events + 1'b1;
                $display("[TB] Backpressure event at time %0t", $time);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Backpressure event at time %0t", $time);
            end
            // Account transactions
            if (valid_in) begin
                if (ready_gated_in)
                    transactions_accepted <= transactions_accepted + 1'b1;
                else
                    transactions_stalled  <= transactions_stalled + 1'b1;
            end
        end
    end
endmodule

/*
 * SCuM-V Controller Integration Testbench with TileLink Echo & Inspection
 * 
 * This testbench instantiates the complete a7top module and tests the STL
 * functionality by reading UART byte streams generated by tl_host_sim.py
 * and feeding them through a UART transmitter to simulate real host communication.
 * 
 * TileLink Echo Architecture:
 * - TL_OUT → GenericDeserializer (packet inspection) → GenericSerializer → TL_IN
 * - Provides realistic echo behavior with proper serialization/deserialization timing
 * - Captures complete TileLink packets for validation and debugging
 * 
 * Test flow:
 * 1. Read test vector file generated by tl_host_sim.py
 * 2. Feed bytes through UART transmitter to generate proper UART timing
 * 3. Connect UART output to a7top UART input
 * 4. TileLink packets sent via TL_OUT are echoed back via TL_IN
 * 5. GenericDeserializer inspects packets and displays all fields
 * 6. Comprehensive validation with content-based assertions
 * 7. Capture and verify UART response packets
 * 
 * Validation Features:
 * - Echo functionality: Commands are properly echoed back
 * - Packet inspection: Deserialized packets show exactly what was transmitted
 * - Content validation: Assertions verify packet field validity
 * - Pass/fail criteria: UART responses + TileLink packets + assertion results
 * 
 * Usage with Vivado:
 * 1. Generate test vectors: python tl_host_sim.py --generate-test-vectors -o sim_input.bin
 * 2. Run simulation with: sim:/scumv_controller_integration_tb
 */

// Dual logging implemented explicitly at each callsite using $display and $fdisplay

module scumv_controller_integration_tb();

    // Test parameters
    parameter CLOCK_FREQ = 100_000_000;  // 100 MHz system clock
    parameter BAUD_RATE = 2_000_000;     // UART baud rate
    parameter TEST_VECTOR_FILE = "C:/Projects/Repositories/scum-v-bringup/hw/scumv-controller/sim/stl_flash_stress_4096pkts.bin";  // Input file from tl_host_sim.py
    parameter MAX_BYTES = 1048576;       // Maximum test vector size (1 MiB)
    parameter TIMEOUT_CYCLES = 5000000;  // Timeout for waiting operations
    parameter STOP_ON_FAIL   = 1;        // Pause simulation on first assertion failure

    // STL batching parameters to mimic tl_host.py batched streaming
    parameter PACKET_LEN_STL = 20;            // 4-byte "stl+" prefix + 16-byte TL payload
    parameter PACKETS_PER_BATCH = 64;         // Number of STL packets per batch
    parameter INTER_BYTE_GAP_CYCLES = 0;      // Extra gaps beyond UART stop bit (keep 0)
    parameter BATCH_DELAY_TL_CYCLES = 16;      // TL clock cycles to wait between batches

    // SerDes backpressure modeling parameters
    parameter SERDES_BACKPRESSURE_ENABLE = 1;  // Enable/disable backpressure modeling
    parameter SERDES_PATTERN_LEN = 9;          // Length of the backpressure pattern
    
    // Clock and reset
    reg clk;
    reg reset_n;
    wire reset = ~reset_n;

    // Log file descriptor for mirroring $display output to a file
    integer tb_log_fd;
    
    // Test control
    reg [7:0] test_vectors [0:MAX_BYTES-1];  // Test vector memory
    integer test_vector_size;                 // Actual size of loaded vectors
    integer current_byte;                     // Current byte being sent
    reg test_active;                          // Test is running
    reg [31:0] timeout_counter;               // Timeout counter
    integer stl_packet_count_total;           // Count of STL packets detected in input
    integer packet_offsets [0:MAX_BYTES-1];   // Byte offsets for each detected STL packet
    
    // UART stimulus generation
    reg [7:0] uart_tx_data;
    reg uart_tx_valid;
    wire uart_tx_ready;
    wire uart_tx_serial;
    
    // UART response capture
    wire [7:0] uart_rx_data;
    wire uart_rx_valid;
    reg uart_rx_ready;
    wire uart_rx_serial;
    reg [7:0] response_buffer [0:255];       // Response capture buffer
    integer response_count;                   // Number of response bytes received
    
    // Device under test (DUT) - a7top module
    wire [3:0] led;
    
    // SerialTL interface - now with loopback and inspection
    reg tl_clk;
    wire tl_in_valid;
    wire tl_in_ready;
    wire tl_in_data;
    wire tl_out_valid;
    wire tl_out_ready;
    wire tl_out_data;
    
    // TileLink packet inspection signals
    wire tl_inspector_ready;
    wire tl_inspector_valid;
    wire [2:0] tl_inspector_chanId;
    wire [2:0] tl_inspector_opcode;
    wire [2:0] tl_inspector_param;
    wire [7:0] tl_inspector_size;
    wire [7:0] tl_inspector_source;
    wire [63:0] tl_inspector_address;
    wire [63:0] tl_inspector_data;
    wire tl_inspector_corrupt;
    wire [8:0] tl_inspector_union;
    // Simple ready/valid handshake between deserializer (producer) and serializer (consumer)
    wire ser_in_ready; // serializer input readiness fed back to deserializer

    // SerDes backpressure modeling: patterns and intermediate signals
    reg [8:0] tl_in_ready_pattern;
    reg [8:0] tl_out_ready_pattern;
    wire [3:0] tl_in_ready_cnt_idx;
    wire [3:0] tl_out_ready_cnt_idx;
    wire tl_in_ready_gated;      // Gated ready seen by serializer output
    wire tl_out_ready_gated;     // Gated ready seen by DUT on TL_OUT
    wire ser_to_dut_valid;       // Serializer to DUT valid
    wire ser_to_dut_ready;       // DUT actual ready (raw)
    wire dut_to_deser_ready;     // Deserializer actual ready (raw)

    // Backpressure counters (exposed for reporting)
    wire [31:0] tl_in_backpressure_events;
    wire [31:0] tl_out_backpressure_events;
    wire [31:0] tl_in_transactions_accepted;
    wire [31:0] tl_in_transactions_stalled;
    wire [31:0] tl_out_transactions_accepted;
    wire [31:0] tl_out_transactions_stalled;
    
    // Mock ASC interface
    wire scan_clk, scan_en, scan_in, scan_reset;

    // Initialize backpressure patterns
    initial begin
        tl_in_ready_pattern  = 9'b111111110;   // 8 cycles accept, 1 cycle backpressure
        tl_out_ready_pattern = 9'b111111110;   // 8 cycles accept, 1 cycle backpressure
    end
    
    // TileLink packet inspector (deserializer for monitoring)
    GenericDeserializer tl_inspector (
        .clock(tl_clk),
        .reset(reset),
        .io_in_ready(tl_inspector_ready),    // Deserializer raw ready
        .io_in_valid(tl_out_valid),          // Direct from DUT TL_OUT
        .io_in_bits(tl_out_data),            // Input from DUT TL_OUT
        .io_out_ready(ser_in_ready),         // Serializer's actual ready signal
        .io_out_valid(tl_inspector_valid),
        .io_out_bits_chanId(tl_inspector_chanId),
        .io_out_bits_opcode(tl_inspector_opcode),
        .io_out_bits_param(tl_inspector_param),
        .io_out_bits_size(tl_inspector_size),
        .io_out_bits_source(tl_inspector_source),
        .io_out_bits_address(tl_inspector_address),
        .io_out_bits_data(tl_inspector_data),
        .io_out_bits_corrupt(tl_inspector_corrupt),
        .io_out_bits_union(tl_inspector_union)
    );
    
    // TileLink echo serializer (re-serializes packets back to TL_IN)
    GenericSerializer tl_echo_serializer (
        .clock(tl_clk),
        .reset(reset),
        .io_in_ready(ser_in_ready),              // Feed back to deserializer for proper handshake
        .io_in_valid(tl_inspector_valid),        // Input from deserializer
        .io_in_bits_chanId(tl_inspector_chanId),
        .io_in_bits_opcode(tl_inspector_opcode),
        .io_in_bits_param(tl_inspector_param),
        .io_in_bits_size(tl_inspector_size),
        .io_in_bits_source(tl_inspector_source),
        .io_in_bits_address(tl_inspector_address),
        .io_in_bits_data(tl_inspector_data),
        .io_in_bits_corrupt(tl_inspector_corrupt),
        .io_in_bits_union(tl_inspector_union),
        .io_in_bits_last(1'b1),                 // Always last bit for single packets
        .io_out_ready(tl_in_ready_gated),       // Gated ready towards serializer output
        .io_out_valid(ser_to_dut_valid),        // Serializer's valid output
        .io_out_bits(tl_in_data)                 // Output to DUT TL_IN
    );
    
    // Ready gating and counters: TL_IN path (Serializer → DUT)
    assign ser_to_dut_ready = tl_in_ready;  // DUT actual ready (raw)
    rv_ready_gate #(.PATTERN_LEN(SERDES_PATTERN_LEN)) gate_tl_in (
        .clock(tl_clk),
        .reset(reset),
        .enable(SERDES_BACKPRESSURE_ENABLE),
        .pattern(tl_in_ready_pattern),
        .valid_in(ser_to_dut_valid),
        .raw_ready_in(ser_to_dut_ready),
        .index(tl_in_ready_cnt_idx),
        .ready_gated_out(tl_in_ready_gated)
    );
    rv_bp_counters cnt_tl_in (
        .clock(tl_clk),
        .reset(reset),
        .enable(SERDES_BACKPRESSURE_ENABLE),
        .valid_in(ser_to_dut_valid),
        .raw_ready_in(ser_to_dut_ready),
        .ready_gated_in(tl_in_ready_gated),
        .tb_log_fd(tb_log_fd),
        .backpressure_events(tl_in_backpressure_events),
        .transactions_accepted(tl_in_transactions_accepted),
        .transactions_stalled(tl_in_transactions_stalled)
    );

    // Ready gating and counters: TL_OUT path (DUT → Deserializer)
    assign dut_to_deser_ready = tl_inspector_ready; // Deserializer actual raw ready
    rv_ready_gate #(.PATTERN_LEN(SERDES_PATTERN_LEN)) gate_tl_out (
        .clock(tl_clk),
        .reset(reset),
        .enable(SERDES_BACKPRESSURE_ENABLE),
        .pattern(tl_out_ready_pattern),
        .valid_in(tl_out_valid),
        .raw_ready_in(dut_to_deser_ready),
        .index(tl_out_ready_cnt_idx),
        .ready_gated_out(tl_out_ready_gated)
    );
    rv_bp_counters cnt_tl_out (
        .clock(tl_clk),
        .reset(reset),
        .enable(SERDES_BACKPRESSURE_ENABLE),
        .valid_in(tl_out_valid),
        .raw_ready_in(dut_to_deser_ready),
        .ready_gated_in(tl_out_ready_gated),
        .tb_log_fd(tb_log_fd),
        .backpressure_events(tl_out_backpressure_events),
        .transactions_accepted(tl_out_transactions_accepted),
        .transactions_stalled(tl_out_transactions_stalled)
    );

    // Final connections to DUT with gated ready
    assign tl_in_valid = ser_to_dut_valid;       // Direct connection (no masking)
    assign tl_out_ready = tl_out_ready_gated;    // What DUT sees on TL_OUT ready
    // Valid is not gated into deserializer; only ready is patterned

    // Test validation variables
    integer packets_sent_count;
    integer packets_received_count;
    integer assertion_failures;
    integer prev_assertion_failures;
    reg test_passed;
    integer expected_pkt_index;               // Index into expected STL packets for comparisons
    // Expected-packet scratch registers (declared at module scope for Verilog-2001 compatibility)
    integer base_idx;
    reg [7:0] chanid_b, opcode_packed_b, size_b, union_b;
    reg [31:0] addr32_le;
    reg [63:0] data64_le;
    reg [2:0] exp_chanid, exp_opcode, exp_param;
    reg [7:0] exp_size, exp_source;
    reg [63:0] exp_addr64, exp_data64;
    reg       exp_corrupt;
    reg [8:0] exp_union9;
    
    // UART stimulus generator (transmitter to feed data to DUT)
    uart #(
        .CLOCK_FREQ(CLOCK_FREQ),
        .BAUD_RATE(BAUD_RATE)
    ) uart_stimulus (
        .clk(clk),
        .reset(reset),
        .data_in(uart_tx_data),
        .data_in_valid(uart_tx_valid),
        .data_in_ready(uart_tx_ready),
        .data_out(),           // Not used for stimulus
        .data_out_valid(),     // Not used for stimulus  
        .data_out_ready(1'b0), // Not used for stimulus
        .serial_in(1'b1),      // Idle state
        .serial_out(uart_tx_serial)
    );
    
    // UART response capture (receiver to capture responses from DUT)
    uart #(
        .CLOCK_FREQ(CLOCK_FREQ),
        .BAUD_RATE(BAUD_RATE)
    ) uart_capture (
        .clk(clk),
        .reset(reset),
        .data_in(8'h00),       // Not used for capture
        .data_in_valid(1'b0),  // Not used for capture
        .data_in_ready(),      // Not used for capture
        .data_out(uart_rx_data),
        .data_out_valid(uart_rx_valid),
        .data_out_ready(uart_rx_ready),
        .serial_in(uart_rx_serial),  // Connected to DUT UART output
        .serial_out()          // Not used for capture
    );
    
    // Device Under Test - SCuM-V Controller
    a7top dut (
        .CLK100MHZ(clk),
        .RESET(reset_n),  // a7top expects active-high reset, reset_n is active-low
        .BUTTON_0(1'b1),   // Button not pressed (active-low)
        .led(led),
        
        // UART interface
        .UART_TXD_IN(uart_tx_serial),      // Input to FPGA from our stimulus generator
        .UART_RXD_IN(uart_rx_serial),      // Output from FPGA to our response capture
        
        // SerialTL interface (mocked)
        .TL_CLK(tl_clk),
        .TL_IN_VALID(tl_in_valid),
        .TL_IN_READY(tl_in_ready),
        .TL_IN_DATA(tl_in_data),
        .TL_OUT_VALID(tl_out_valid),
        .TL_OUT_READY(tl_out_ready),
        .TL_OUT_DATA(tl_out_data),
        
        // ASC interface (not used in this test) 
        .SCAN_CLK(scan_clk),
        .SCAN_EN(scan_en),
        .SCAN_IN(scan_in),
        .SCAN_RESET(scan_reset),
        .CHIP_RESET()  // Not connected in this test
    );
    
    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // 100 MHz clock (10ns period)
    end
    
    // TileLink clock generation (mock - 50 kHz)
    initial begin
        tl_clk = 0;
        forever #1000 tl_clk = ~tl_clk;  // 500 kHz TL clock (period = 2 us, half-period = 1 us = 1000 ns)
    end
    
    // Main test procedure
    initial begin
        // Open log file early so all subsequent messages are mirrored to file as well
        tb_log_fd = $fopen("scumv_controller_integration_tb.log", "w");
        $display("[TB] Starting SCuM-V Controller Integration Test");
        if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Starting SCuM-V Controller Integration Test");
        $display("[TB] Clock Freq: %0d Hz, BAUD Rate: %0d", CLOCK_FREQ, BAUD_RATE);
        if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Clock Freq: %0d Hz, BAUD Rate: %0d", CLOCK_FREQ, BAUD_RATE);
        
        // Initialize signals
        reset_n = 0;
        uart_tx_data = 8'h00;
        uart_tx_valid = 1'b0;
        uart_rx_ready = 1'b1;  // Always ready to receive responses
        current_byte = 0;
        test_active = 1'b0;
        response_count = 0;
        timeout_counter = 0;
        
        // Initialize test validation variables
        packets_sent_count = 0;
        packets_received_count = 0;
        assertion_failures = 0;
        prev_assertion_failures = 0;
        test_passed = 1'b0;
        expected_pkt_index = 0;
        
        // TileLink interface is now active with loopback connections
        // (no initialization needed - handled by assign statements)
        
        // Load test vectors from file
        load_test_vectors();
        
        // Reset sequence
        $display("[TB] Applying reset...");
        if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Applying reset...");
        #12000;
        reset_n = 1;
        #12000;
        $display("[TB] Reset released, starting test sequence");
        if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Reset released, starting test sequence");
        
        // Wait for system to settle
        #1000;
        
        // Start test sequence
        test_active = 1'b1;
        send_test_vectors();
        
        // Wait for all responses or timeout
        wait_for_responses();
        
        // Analyze results
        analyze_results();
        
        $display("[TB] Test completed");
        if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Test completed");
        if (tb_log_fd) $fclose(tb_log_fd);
        $finish;
    end

    // Optional: pause simulation on the first assertion failure to aid debugging
    always @(posedge tl_clk) begin
        if (STOP_ON_FAIL && (assertion_failures > prev_assertion_failures)) begin
            $display("[TB] STOP_ON_FAIL: Pausing on first assertion failure at time %0t", $time);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] STOP_ON_FAIL: Pausing on first assertion failure at time %0t", $time);
            $stop; // Pause simulation for interactive debug
        end
        prev_assertion_failures <= assertion_failures;
    end

    // Load test vectors from file
    task load_test_vectors;
        integer file_handle, byte_val, i;
        begin
            $display("[TB] Loading test vectors from %s", TEST_VECTOR_FILE);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Loading test vectors from %s", TEST_VECTOR_FILE);
            
            file_handle = $fopen(TEST_VECTOR_FILE, "rb");
            if (file_handle == 0) begin
                $display("[TB] ERROR: Could not open test vector file %s", TEST_VECTOR_FILE);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ERROR: Could not open test vector file %s", TEST_VECTOR_FILE);
                $display("[TB] Please run: python tl_host_sim.py --generate-test-vectors -o %s", TEST_VECTOR_FILE);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Please run: python tl_host_sim.py --generate-test-vectors -o %s", TEST_VECTOR_FILE);
                $finish;
            end
            
            test_vector_size = 0;
            for (i = 0; i < MAX_BYTES; i = i + 1) begin
                byte_val = $fgetc(file_handle);
                if (byte_val == -1) begin
                    i = MAX_BYTES;  // Exit loop on EOF
                end else begin
                    test_vectors[i] = byte_val[7:0];
                    test_vector_size = test_vector_size + 1;
                end
            end
            
            $fclose(file_handle);
            $display("[TB] Loaded %0d bytes from test vector file", test_vector_size);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Loaded %0d bytes from test vector file", test_vector_size);
            
            // Display first few bytes for debugging
            $write("[TB] First 16 bytes: ");
            for (i = 0; i < 16 && i < test_vector_size; i = i + 1) begin
                $write("%02X ", test_vectors[i]);
            end
            $write("\n");
        end
    endtask
    
    // Count STL packets by scanning for "stl+" prefix every PACKET_LEN_STL bytes
    task count_stl_packets;
        integer i, j, preview_end, base0;
        begin
            stl_packet_count_total = 0;
            i = 0;
            while (i + 3 < test_vector_size) begin
                if (test_vectors[i]   == 8'h73 && // 's'
                    test_vectors[i+1] == 8'h74 && // 't'
                    test_vectors[i+2] == 8'h6C && // 'l'
                    test_vectors[i+3] == 8'h2B)   // '+'
                begin
                    packet_offsets[stl_packet_count_total] = i;
                    stl_packet_count_total = stl_packet_count_total + 1;
                    i = i + PACKET_LEN_STL;
                end else begin
                    // Advance by one to allow misalignment detection
                    i = i + 1;
                end
            end
            $display("[TB] Detected %0d STL packets (PACKET_LEN_STL=%0d)", stl_packet_count_total, PACKET_LEN_STL);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Detected %0d STL packets (PACKET_LEN_STL=%0d)", stl_packet_count_total, PACKET_LEN_STL);
            if (stl_packet_count_total > 0) begin
                base0 = packet_offsets[0];
                preview_end = (base0 + 8 <= test_vector_size) ? base0 + 8 : test_vector_size;
                $write("[TB] First packet bytes at offset %0d: ", base0);
                for (j = base0; j < preview_end; j = j + 1) $write("%02X ", test_vectors[j]);
                $write("\n");
            end
        end
    endtask
    
    // Send a batch of STL packets continuously over UART (mimics tl_host batched streaming)
    task send_stl_batch(input integer start_packet_idx, input integer num_packets);
        integer pkt, byte_idx, base_idx, tl_pause_cnt;
        begin
            for (pkt = 0; pkt < num_packets; pkt = pkt + 1) begin
                base_idx = packet_offsets[start_packet_idx + pkt];
                // Send one full 20-byte STL command: "stl+" + 16B TL payload
                for (byte_idx = 0; byte_idx < PACKET_LEN_STL; byte_idx = byte_idx + 1) begin
                    // Ensure transmitter is ready before presenting the byte
                    wait_for_uart_ready();
                    uart_tx_data  = test_vectors[base_idx + byte_idx];
                    uart_tx_valid = 1'b1;
                    @(posedge clk);
                    // Confirm transmitter has started (ready dropped), then release VALID
                    wait (!uart_tx_ready);
                    uart_tx_valid = 1'b0;
                    // Wait until transmitter finishes current byte (ready high again)
                    wait (uart_tx_ready);
                    // Optional minimal gap between bytes (keep 0 to stress DUT)
                    repeat(INTER_BYTE_GAP_CYCLES) @(posedge clk);
                end
                packets_sent_count = packets_sent_count + 1;
            $display("[TB] Sent STL packet #%0d (byte range %0d..%0d)",
                         start_packet_idx + pkt,
                         base_idx,
                         base_idx + PACKET_LEN_STL - 1);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Sent STL packet #%0d (byte range %0d..%0d)",
                         start_packet_idx + pkt,
                         base_idx,
                         base_idx + PACKET_LEN_STL - 1);
            end
            // Optional pause between batches to emulate host think time
            if (BATCH_DELAY_TL_CYCLES > 0) begin
                for (tl_pause_cnt = 0; tl_pause_cnt < BATCH_DELAY_TL_CYCLES; tl_pause_cnt = tl_pause_cnt + 1)
                    @(posedge tl_clk);
            end
        end
    endtask

    // Send test vectors as STL packets in batches (no artificial per-byte delays)
    task send_test_vectors;
        integer total_batches, b, remaining, count_this_batch, start_pkt;
        begin
            $display("[TB] Preparing to send STL packets in batches of %0d", PACKETS_PER_BATCH);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Preparing to send STL packets in batches of %0d", PACKETS_PER_BATCH);
            count_stl_packets();

            total_batches = (stl_packet_count_total + PACKETS_PER_BATCH - 1) / PACKETS_PER_BATCH;
            for (b = 0; b < total_batches; b = b + 1) begin
                start_pkt = b * PACKETS_PER_BATCH;
                remaining = stl_packet_count_total - start_pkt;
                count_this_batch = (remaining > PACKETS_PER_BATCH) ? PACKETS_PER_BATCH : remaining;
                $display("[TB] Sending batch %0d/%0d: %0d packets (start index %0d)",
                         b+1, total_batches, count_this_batch, start_pkt);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Sending batch %0d/%0d: %0d packets (start index %0d)",
                         b+1, total_batches, count_this_batch, start_pkt);
                send_stl_batch(start_pkt, count_this_batch);
            end
            $display("[TB] All STL packets sent: %0d", stl_packet_count_total);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] All STL packets sent: %0d", stl_packet_count_total);
        end
    endtask
    
    // Wait for UART transmitter to be ready
    task wait_for_uart_ready;
        begin
            timeout_counter = 0;
            while (!uart_tx_ready && timeout_counter < TIMEOUT_CYCLES) begin
                @(posedge clk);
                timeout_counter = timeout_counter + 1;
            end
            
            if (timeout_counter >= TIMEOUT_CYCLES) begin
            $display("[TB] ERROR: Timeout waiting for UART TX ready");
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ERROR: Timeout waiting for UART TX ready");
                $finish;
            end
        end
    endtask
    
    // Wait for responses from DUT
    task wait_for_responses;
        integer expected_bytes;
        begin
            expected_bytes = packets_sent_count * 16; // 16 bytes per STL response
            $display("[TB] Waiting for %0d response bytes (for %0d packets)", expected_bytes, packets_sent_count);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Waiting for %0d response bytes (for %0d packets)", expected_bytes, packets_sent_count);
            timeout_counter = 0;

            while ((response_count < expected_bytes) && (timeout_counter < TIMEOUT_CYCLES)) begin
                @(posedge clk);
                timeout_counter = timeout_counter + 1;
            end

            if (response_count < expected_bytes) begin
                $display("[TB] ERROR: Expected %0d response bytes, got %0d", expected_bytes, response_count);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ERROR: Expected %0d response bytes, got %0d", expected_bytes, response_count);
                assertion_failures = assertion_failures + 1;
            end else begin
                $display("[TB] Collected expected %0d response bytes", response_count);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Collected expected %0d response bytes", response_count);
            end
        end
    endtask
    
    // Analyze test results
    task analyze_results;
        integer i;
        begin
            $display("[TB] ========== TEST RESULTS ==========");
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ========== TEST RESULTS ==========");
            $display("[TB] Test vectors sent: %0d bytes", test_vector_size);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Test vectors sent: %0d bytes", test_vector_size);
            $display("[TB] Response bytes received: %0d", response_count);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Response bytes received: %0d", response_count);
            
            if (response_count > 0) begin
                $write("[TB] Response bytes: ");
                for (i = 0; i < response_count && i < 32; i = i + 1) begin
                    $write("%02X ", response_buffer[i]);
                end
                if (response_count > 32) $write("... (truncated)");
                $write("\n");
            end
            
            // TileLink packet validation results
            $display("[TB] TileLink packets received: %0d", packets_received_count);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] TileLink packets received: %0d", packets_received_count);
            $display("[TB] Assertion failures: %0d", assertion_failures);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Assertion failures: %0d", assertion_failures);
            
            // Check LED status
            $display("[TB] Final LED status: %b", led);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Final LED status: %b", led);
            $display("[TB] LED[0] (n_reset): %b", led[0]);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] LED[0] (n_reset): %b", led[0]); 
            $display("[TB] LED[1] (ASC active): %b", led[1]); 
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] LED[1] (ASC active): %b", led[1]); 
            $display("[TB] LED[2] (STL active): %b", led[2]);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] LED[2] (STL active): %b", led[2]);
            $display("[TB] LED[3] (TL_IN_VALID): %b", led[3]);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] LED[3] (TL_IN_VALID): %b", led[3]);
            
            // Backpressure statistics
            if (SERDES_BACKPRESSURE_ENABLE) begin
                $display("[TB] ========== BACKPRESSURE STATISTICS ==========");
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ========== BACKPRESSURE STATISTICS ==========");
                
                $display("[TB] TL_IN Path (Serializer → DUT):");
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] TL_IN Path (Serializer → DUT):");
                $display("[TB]   Pattern: %b", tl_in_ready_pattern);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB]   Pattern: %b", tl_in_ready_pattern);
                $display("[TB]   Transactions accepted: %0d", tl_in_transactions_accepted);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB]   Transactions accepted: %0d", tl_in_transactions_accepted);
                $display("[TB]   Transactions stalled: %0d", tl_in_transactions_stalled);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB]   Transactions stalled: %0d", tl_in_transactions_stalled);
                $display("[TB]   Backpressure events: %0d", tl_in_backpressure_events);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB]   Backpressure events: %0d", tl_in_backpressure_events);
                
                $display("[TB] TL_OUT Path (DUT → Deserializer):");
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] TL_OUT Path (DUT → Deserializer):");
                $display("[TB]   Pattern: %b", tl_out_ready_pattern);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB]   Pattern: %b", tl_out_ready_pattern);
                $display("[TB]   Transactions accepted: %0d", tl_out_transactions_accepted);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB]   Transactions accepted: %0d", tl_out_transactions_accepted);
                $display("[TB]   Transactions stalled: %0d", tl_out_transactions_stalled);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB]   Transactions stalled: %0d", tl_out_transactions_stalled);
                $display("[TB]   Backpressure events: %0d", tl_out_backpressure_events);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB]   Backpressure events: %0d", tl_out_backpressure_events);
                
                // Calculate effective throughput
                if (tl_in_transactions_accepted + tl_in_transactions_stalled > 0) begin
                    $display("[TB]   TL_IN Throughput: %0.1f%%", 
                        100.0 * tl_in_transactions_accepted / 
                        (tl_in_transactions_accepted + tl_in_transactions_stalled));
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB]   TL_IN Throughput: %0.1f%%", 
                        100.0 * tl_in_transactions_accepted / 
                        (tl_in_transactions_accepted + tl_in_transactions_stalled));
                end
                if (tl_out_transactions_accepted + tl_out_transactions_stalled > 0) begin
                    $display("[TB]   TL_OUT Throughput: %0.1f%%", 
                        100.0 * tl_out_transactions_accepted / 
                        (tl_out_transactions_accepted + tl_out_transactions_stalled));
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB]   TL_OUT Throughput: %0.1f%%", 
                        100.0 * tl_out_transactions_accepted / 
                        (tl_out_transactions_accepted + tl_out_transactions_stalled));
                end
            end
            
            // Comprehensive pass/fail criteria
            test_passed = 1'b1;  // Start with pass assumption
            
            if (response_count == 0) begin
                $display("[TB] FAIL: No UART response data received");
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] FAIL: No UART response data received");
                test_passed = 1'b0;
            end else begin
                $display("[TB] PASS: Received %0d UART response bytes", response_count);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] PASS: Received %0d UART response bytes", response_count);
            end
            
            if (packets_received_count == 0) begin
                $display("[TB] FAIL: No TileLink packets captured");
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] FAIL: No TileLink packets captured");
                test_passed = 1'b0;
            end else begin
                $display("[TB] PASS: Captured %0d TileLink packets", packets_received_count);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] PASS: Captured %0d TileLink packets", packets_received_count);
            end
            
            if (assertion_failures > 0) begin
                $display("[TB] FAIL: %0d assertion failures detected", assertion_failures);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] FAIL: %0d assertion failures detected", assertion_failures);
                test_passed = 1'b0;
            end else begin
                $display("[TB] PASS: No assertion failures");
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] PASS: No assertion failures");
            end
            
            // Final test result
            if (test_passed) begin
                $display("[TB] OVERALL RESULT: PASS - Echo functionality working correctly");
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] OVERALL RESULT: PASS - Echo functionality working correctly");
            end else begin
                $display("[TB] OVERALL RESULT: FAIL - Test validation failed");
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] OVERALL RESULT: FAIL - Test validation failed");
            end
            
            $display("[TB] ===================================");
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ===================================");
        end
    endtask
    
    // Response capture process
    always @(posedge clk) begin
        if (reset) begin
            response_count <= 0;
        end else if (uart_rx_valid && uart_rx_ready) begin
            if (response_count < 256) begin
                response_buffer[response_count] <= uart_rx_data;
                response_count <= response_count + 1;
                $display("[TB] Captured response byte %0d: 0x%02X", response_count, uart_rx_data);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Captured response byte %0d: 0x%02X", response_count, uart_rx_data);
            end
        end
    end
    
    // Monitor and validate deserialized TileLink packets
    always @(posedge tl_clk) begin
        if (tl_inspector_valid) begin
            packets_received_count = packets_received_count + 1;
            
            $display("[TB] ========== TILELINK PACKET CAPTURED ==========");
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ========== TILELINK PACKET CAPTURED ==========");
            $display("[TB] Packet #%0d", packets_received_count);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Packet #%0d", packets_received_count);
            $display("[TB] Channel ID: 0x%01X", tl_inspector_chanId);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Channel ID: 0x%01X", tl_inspector_chanId);
            $display("[TB] Opcode:     0x%01X (%s)", tl_inspector_opcode, 
                     tl_inspector_opcode == 3'h0 ? "PutFullData" :
                     tl_inspector_opcode == 3'h1 ? "PutPartialData" :
                     tl_inspector_opcode == 3'h4 ? "Get" :
                     tl_inspector_opcode == 3'h0 ? "AccessAck" :
                     tl_inspector_opcode == 3'h1 ? "AccessAckData" : "Unknown");
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Opcode:     0x%01X (%s)", tl_inspector_opcode, 
                       tl_inspector_opcode == 3'h0 ? "PutFullData" :
                       tl_inspector_opcode == 3'h1 ? "PutPartialData" :
                       tl_inspector_opcode == 3'h4 ? "Get" :
                       tl_inspector_opcode == 3'h0 ? "AccessAck" :
                       tl_inspector_opcode == 3'h1 ? "AccessAckData" : "Unknown");
            $display("[TB] Param:      0x%01X", tl_inspector_param);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Param:      0x%01X", tl_inspector_param);
            $display("[TB] Size:       0x%02X (%0d bytes)", tl_inspector_size, 1 << tl_inspector_size);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Size:       0x%02X (%0d bytes)", tl_inspector_size, 1 << tl_inspector_size);
            $display("[TB] Source:     0x%02X", tl_inspector_source);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Source:     0x%02X", tl_inspector_source);
            $display("[TB] Address:    0x%016X", tl_inspector_address);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Address:    0x%016X", tl_inspector_address);
            $display("[TB] Data:       0x%016X", tl_inspector_data);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Data:       0x%016X", tl_inspector_data);
            $display("[TB] Corrupt:    %b", tl_inspector_corrupt);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Corrupt:    %b", tl_inspector_corrupt);
            $display("[TB] Union:      0x%03X", tl_inspector_union);
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] Union:      0x%03X", tl_inspector_union);
            $display("[TB] =============================================");
            if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] =============================================");
            
            // Basic packet validation assertions (content only, not timing)
            if (tl_inspector_size > 8'h06) begin
                $error("[TB] ASSERTION FAILED: Invalid packet size: 0x%02X (max 0x06)", tl_inspector_size);
                assertion_failures = assertion_failures + 1;
            end
            
            if (tl_inspector_chanId > 3'h2) begin
                $error("[TB] ASSERTION FAILED: Invalid channel ID: 0x%01X (max 0x2)", tl_inspector_chanId);
                assertion_failures = assertion_failures + 1;
            end
            
            if (tl_inspector_opcode > 3'h6) begin
                $error("[TB] ASSERTION FAILED: Invalid opcode: 0x%01X (max 0x6)", tl_inspector_opcode);
                assertion_failures = assertion_failures + 1;
            end

            // Compare deserialized packet against what was sent in the UART STL vector
            // Reconstruct expected fields directly from test_vectors using packet_offsets[]
            // STL packet format: 'stl+' (4B) + 16B TL payload packed as <BBBBLQ>
            //   Byte 0: chanid (3 LSBs used)
            //   Byte 1: opcode_packed = {corrupt[7], param[6:4], 1'b0, opcode[2:0]}
            //   Byte 2: size
            //   Byte 3: union_field (mask for Ch A, denied for Ch D)
            //   Bytes 4..7: address (LE, 32-bit)
            //   Bytes 8..15: data (LE, 64-bit)
            if (expected_pkt_index < stl_packet_count_total) begin
                base_idx = packet_offsets[expected_pkt_index] + 4; // skip 'stl+'
                chanid_b         = test_vectors[base_idx + 0];
                opcode_packed_b  = test_vectors[base_idx + 1];
                size_b           = test_vectors[base_idx + 2];
                union_b          = test_vectors[base_idx + 3];
                addr32_le        = { test_vectors[base_idx + 7], test_vectors[base_idx + 6],
                                      test_vectors[base_idx + 5], test_vectors[base_idx + 4] };
                data64_le        = { test_vectors[base_idx + 15], test_vectors[base_idx + 14],
                                      test_vectors[base_idx + 13], test_vectors[base_idx + 12],
                                      test_vectors[base_idx + 11], test_vectors[base_idx + 10],
                                      test_vectors[base_idx + 9],  test_vectors[base_idx + 8] };

                exp_chanid  = chanid_b[2:0];
                exp_opcode  = opcode_packed_b[2:0];
                exp_param   = opcode_packed_b[6:4];
                exp_corrupt = opcode_packed_b[7];
                exp_size    = size_b;
                exp_source  = 8'h00; // host transactions default source
                exp_union9  = {1'b0, union_b}; // zero-extend to 9 bits
                exp_addr64  = {32'h0, addr32_le};
                exp_data64  = data64_le;

                // Field-by-field comparisons
                if (tl_inspector_chanId !== exp_chanid) begin
                    $error("[TB] ASSERTION FAILED: Packet #%0d chanId mismatch: got 0x%0X expected 0x%0X", expected_pkt_index+1, tl_inspector_chanId, exp_chanid);
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ASSERTION FAILED: Packet #%0d chanId mismatch: got 0x%0X expected 0x%0X", expected_pkt_index+1, tl_inspector_chanId, exp_chanid);
                    assertion_failures = assertion_failures + 1;
                end
                if (tl_inspector_opcode !== exp_opcode) begin
                    $error("[TB] ASSERTION FAILED: Packet #%0d opcode mismatch: got 0x%0X expected 0x%0X", expected_pkt_index+1, tl_inspector_opcode, exp_opcode);
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ASSERTION FAILED: Packet #%0d opcode mismatch: got 0x%0X expected 0x%0X", expected_pkt_index+1, tl_inspector_opcode, exp_opcode);
                    assertion_failures = assertion_failures + 1;
                end
                if (tl_inspector_param !== exp_param) begin
                    $error("[TB] ASSERTION FAILED: Packet #%0d param mismatch: got 0x%0X expected 0x%0X", expected_pkt_index+1, tl_inspector_param, exp_param);
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ASSERTION FAILED: Packet #%0d param mismatch: got 0x%0X expected 0x%0X", expected_pkt_index+1, tl_inspector_param, exp_param);
                    assertion_failures = assertion_failures + 1;
                end
                if (tl_inspector_size !== exp_size) begin
                    $error("[TB] ASSERTION FAILED: Packet #%0d size mismatch: got 0x%0X expected 0x%0X", expected_pkt_index+1, tl_inspector_size, exp_size);
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ASSERTION FAILED: Packet #%0d size mismatch: got 0x%0X expected 0x%0X", expected_pkt_index+1, tl_inspector_size, exp_size);
                    assertion_failures = assertion_failures + 1;
                end
                if (tl_inspector_source !== exp_source) begin
                    $error("[TB] ASSERTION FAILED: Packet #%0d source mismatch: got 0x%0X expected 0x%0X", expected_pkt_index+1, tl_inspector_source, exp_source);
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ASSERTION FAILED: Packet #%0d source mismatch: got 0x%0X expected 0x%0X", expected_pkt_index+1, tl_inspector_source, exp_source);
                    assertion_failures = assertion_failures + 1;
                end
                if (tl_inspector_address !== exp_addr64) begin
                    $error("[TB] ASSERTION FAILED: Packet #%0d address mismatch: got 0x%016X expected 0x%016X", expected_pkt_index+1, tl_inspector_address, exp_addr64);
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ASSERTION FAILED: Packet #%0d address mismatch: got 0x%016X expected 0x%016X", expected_pkt_index+1, tl_inspector_address, exp_addr64);
                    assertion_failures = assertion_failures + 1;
                end
                if (tl_inspector_data !== exp_data64) begin
                    $error("[TB] ASSERTION FAILED: Packet #%0d data mismatch: got 0x%016X expected 0x%016X", expected_pkt_index+1, tl_inspector_data, exp_data64);
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ASSERTION FAILED: Packet #%0d data mismatch: got 0x%016X expected 0x%016X", expected_pkt_index+1, tl_inspector_data, exp_data64);
                    assertion_failures = assertion_failures + 1;
                end
                if (tl_inspector_corrupt !== exp_corrupt) begin
                    $error("[TB] ASSERTION FAILED: Packet #%0d corrupt mismatch: got %0d expected %0d", expected_pkt_index+1, tl_inspector_corrupt, exp_corrupt);
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ASSERTION FAILED: Packet #%0d corrupt mismatch: got %0d expected %0d", expected_pkt_index+1, tl_inspector_corrupt, exp_corrupt);
                    assertion_failures = assertion_failures + 1;
                end
                if (tl_inspector_union !== exp_union9) begin
                    $error("[TB] ASSERTION FAILED: Packet #%0d union mismatch: got 0x%03X expected 0x%03X", expected_pkt_index+1, tl_inspector_union, exp_union9);
                    if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] ASSERTION FAILED: Packet #%0d union mismatch: got 0x%03X expected 0x%03X", expected_pkt_index+1, tl_inspector_union, exp_union9);
                    assertion_failures = assertion_failures + 1;
                end

                expected_pkt_index = expected_pkt_index + 1;
            end else begin
                $display("[TB] WARN: Received more TL packets than STL vectors (%0d > %0d)", expected_pkt_index+1, stl_packet_count_total);
                if (tb_log_fd) $fdisplay(tb_log_fd, "[TB] WARN: Received more TL packets than STL vectors (%0d > %0d)", expected_pkt_index+1, stl_packet_count_total);
                assertion_failures = assertion_failures + 1;
            end
        end
    end
    
    // Monitor for test timeout
    always @(posedge clk) begin
        if (test_active && timeout_counter > TIMEOUT_CYCLES) begin
            $display("[TB] ERROR: Test timeout exceeded");
            $finish;
        end
    end

endmodule
